module core( // modulo de um core
  input clk, // clock
  input resetn, // reset que ativa em zero
  input [31:0] data_in, // dado de entrada
  output reg [31:0] data_out, // dado de saída
  output reg [31:0] address, // endereço de saída
  output reg we // write enable
);

always @(posedge clk) begin
  if (resetn == 1'b0) begin
    address <= 32'h00000000;
  end else begin
    address <= address + 4;
  end
  we = 0;
  data_out = 32'h00000000;
end

endmodule
